--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   20:10:07 03/10/2016
-- Design Name:   
-- Module Name:   C:/Users/Kristian/Documents/Github/Repositories/4. Semester/Mit/DIG/Projects/Portefolje_1/tb_cnt999.vhd
-- Project Name:  Portefolje_1
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: cnt999
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY tb_cnt999 IS
END tb_cnt999;
 
ARCHITECTURE behavior OF tb_cnt999 IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT cnt999
    PORT(
         clk : IN  std_logic;
         clr : IN  std_logic;
         en : IN  std_logic;
         co : OUT  std_logic;
         bcd : OUT  std_logic_vector(3 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal clr : std_logic := '0';
   signal en : std_logic := '1';

 	--Outputs
   signal co : std_logic;
   signal bcd : std_logic_vector(3 downto 0);

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: cnt999 PORT MAP (
          clk => clk,
          clr => clr,
          en => en,
          co => co,
          bcd => bcd
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;
 
      wait for clk_period*100;
		
		clr <= '1';
		
		wait for 50 ns;
		
		clr <= '0';

      -- insert stimulus here 

      wait;
   end process;

END;
